module fiveBitFullAdder(A, B, Ci, Co, S);
  input wire [4:0] A, B;
  input wire Ci;
  output wire [4:0] S;
  output wire Co;
  wire [4:0] C;

  oneBitFullAdder s1(A[0], B[0], Ci, C[0], S[0]);
  oneBitFullAdder s2(A[1], B[1], C[0], C[1], S[1]);
  oneBitFullAdder s3(A[2], B[2], C[1], C[2], S[2]);
  oneBitFullAdder s4(A[3], B[3], C[2], C[3], S[3]);
  oneBitFullAdder s5(A[4], B[4], C[3], C[4], S[4]);

  assign Co = C[4];
endmodule
