library verilog;
use verilog.vl_types.all;
entity fDDNF is
    port(
        x3              : in     vl_logic;
        x2              : in     vl_logic;
        x1              : in     vl_logic;
        \out\           : out    vl_logic
    );
end fDDNF;
